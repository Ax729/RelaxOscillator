magic
tech sky130A
magscale 1 2
timestamp 1761868743
<< nwell >>
rect -2876 -331 -2079 -10
rect -1173 -331 3550 -10
rect -2796 -1474 -2079 -1410
rect -2900 -1642 -2079 -1474
rect -2796 -1731 -2079 -1642
rect -2044 -1731 -1226 -1410
rect -1173 -1731 3308 -1410
<< pwell >>
rect -2661 829 -2311 1011
rect -2859 -571 -2179 -389
rect -1067 -571 3421 -389
rect -2859 -1971 -2179 -1789
rect -1225 -1971 3419 -1789
rect -2659 -3069 -2321 -2887
<< viali >>
rect -2173 1023 -2123 1067
rect -1740 1060 -1700 1100
rect -1585 1023 -1535 1063
rect -2235 -377 -2197 -339
rect -1614 -356 -1570 -312
rect -1201 -377 -1151 -337
rect -78 -377 -28 -327
rect 498 -373 532 -339
rect 1345 -377 1379 -337
rect 2020 -377 2054 -337
rect 2536 -378 2570 -344
rect 3316 -377 3350 -337
rect 4100 -386 4142 -340
rect -1959 -1771 -1925 -1737
rect -1610 -1756 -1562 -1712
rect -1285 -1777 -1235 -1737
rect -76 -1777 -26 -1727
rect 505 -1777 539 -1743
rect 1479 -1777 1513 -1737
rect 1950 -1777 1984 -1737
rect 2519 -1779 2553 -1745
rect 3314 -1777 3348 -1737
rect 4102 -1778 4138 -1738
rect -2352 -2875 -2301 -2831
rect -1748 -2844 -1710 -2808
rect -1511 -2875 -1461 -2835
<< metal1 >>
rect -2591 1385 -2457 1400
rect -2615 1380 -2352 1385
rect -2664 1304 -2352 1380
rect -2664 1184 -2568 1304
rect -2670 1088 -2664 1184
rect -2568 1088 -2562 1184
rect -1760 1100 -1680 1122
rect -2194 1067 -2108 1082
rect -2194 1023 -2173 1067
rect -2123 1023 -2108 1067
rect -1760 1060 -1740 1100
rect -1700 1090 -1680 1100
rect -1598 1090 -1520 1100
rect -1700 1064 -1520 1090
rect -1700 1063 -780 1064
rect -1700 1060 -1585 1063
rect -1760 1058 -1585 1060
rect -1760 1042 -1680 1058
rect -2194 1004 -2108 1023
rect -1598 1023 -1585 1058
rect -1535 1023 -780 1063
rect -1598 1010 -1520 1023
rect -2174 972 -2124 1004
rect -2921 922 -2124 972
rect -3162 786 -2397 856
rect -3162 760 -2463 786
rect -3162 -544 -3066 760
rect -2664 586 -2568 592
rect -2664 0 -2568 490
rect -824 144 -780 1023
rect -834 92 -828 144
rect -776 92 -770 144
rect -2797 -21 -2275 0
rect -969 -21 3269 0
rect -2797 -31 3269 -21
rect -2784 -47 3251 -31
rect -2784 -65 3271 -47
rect -2797 -96 3271 -65
rect -2664 -262 -2568 -96
rect -828 -194 -776 -188
rect -1614 -242 -828 -198
rect -2670 -358 -2664 -262
rect -2568 -358 -2562 -262
rect -1614 -288 -1570 -242
rect -776 -242 -482 -198
rect -828 -252 -776 -246
rect -1638 -312 -1546 -288
rect -2241 -339 -2191 -327
rect -2241 -377 -2235 -339
rect -2197 -377 -2191 -339
rect -2241 -426 -2191 -377
rect -1638 -356 -1614 -312
rect -1570 -356 -1546 -312
rect -1638 -380 -1546 -356
rect -1220 -337 -1130 -316
rect -1220 -377 -1201 -337
rect -1151 -377 -1130 -337
rect -1220 -400 -1130 -377
rect -533 -326 -482 -242
rect -104 -326 -6 -302
rect -533 -327 -6 -326
rect -533 -377 -78 -327
rect -28 -377 -6 -327
rect -2248 -478 -2242 -426
rect -2190 -478 -2184 -426
rect -1199 -442 -1153 -400
rect -533 -429 -482 -377
rect -104 -396 -6 -377
rect 486 -336 544 -333
rect 1322 -336 1406 -324
rect 486 -337 1406 -336
rect 486 -339 1345 -337
rect 486 -373 498 -339
rect 532 -373 1345 -339
rect 486 -377 1345 -373
rect 1379 -377 1406 -337
rect 486 -379 544 -377
rect 1322 -390 1406 -377
rect 2002 -337 2070 -324
rect 2002 -377 2020 -337
rect 2054 -377 2070 -337
rect 2002 -400 2070 -377
rect 2524 -344 2582 -338
rect 2745 -344 2751 -336
rect 2524 -378 2536 -344
rect 2570 -378 2751 -344
rect 2524 -379 2751 -378
rect 2524 -384 2582 -379
rect 2745 -388 2751 -379
rect 2803 -344 2809 -336
rect 3298 -337 3366 -320
rect 3298 -344 3316 -337
rect 2803 -377 3316 -344
rect 3350 -377 3366 -337
rect 2803 -379 3366 -377
rect 2803 -388 2809 -379
rect 3298 -400 3366 -379
rect 4076 -340 4162 -318
rect 4076 -386 4100 -340
rect 4142 -386 4491 -340
rect -533 -435 -481 -429
rect -1202 -448 -1150 -442
rect 2020 -440 2054 -400
rect 4076 -404 4162 -386
rect -533 -493 -481 -487
rect 2011 -446 2063 -440
rect -1202 -506 -1150 -500
rect 2011 -504 2063 -498
rect -3162 -563 -2325 -544
rect -941 -562 3269 -544
rect -3162 -611 -2130 -563
rect -941 -575 3446 -562
rect -898 -609 3446 -575
rect -3162 -640 -2305 -611
rect -921 -615 3446 -609
rect -921 -640 3293 -615
rect -3162 -1945 -3066 -640
rect -1208 -832 -1202 -780
rect -1150 -783 -1144 -780
rect 2284 -783 2290 -780
rect -1150 -829 2290 -783
rect -1150 -832 -1144 -829
rect 2284 -832 2290 -829
rect 2342 -832 2348 -780
rect -2664 -838 -2568 -832
rect -2664 -1400 -2568 -934
rect 2887 -1213 2893 -1208
rect -1960 -1254 2893 -1213
rect -1960 -1292 -1919 -1254
rect 2887 -1260 2893 -1254
rect 2945 -1260 2951 -1208
rect -1972 -1344 -1966 -1292
rect -1914 -1344 -1908 -1292
rect -2801 -1423 3305 -1400
rect -2811 -1468 3322 -1423
rect -2805 -1495 3305 -1468
rect -2664 -1730 -2568 -1495
rect -1285 -1546 -1233 -1540
rect -1967 -1580 -1915 -1574
rect -1967 -1638 -1915 -1632
rect -1285 -1604 -1233 -1598
rect -1962 -1720 -1921 -1638
rect -1634 -1712 -1540 -1690
rect -2670 -1826 -2664 -1730
rect -2568 -1826 -2562 -1730
rect -1976 -1737 -1914 -1720
rect -1976 -1771 -1959 -1737
rect -1925 -1771 -1914 -1737
rect -1976 -1786 -1914 -1771
rect -1634 -1756 -1610 -1712
rect -1562 -1756 -1540 -1712
rect -1285 -1714 -1234 -1604
rect 2504 -1612 2510 -1560
rect 2562 -1612 2568 -1560
rect 2892 -1588 2944 -1582
rect 917 -1658 1984 -1624
rect -1634 -1780 -1540 -1756
rect -1306 -1737 -1218 -1714
rect -94 -1726 -8 -1710
rect -1306 -1777 -1285 -1737
rect -1235 -1777 -1218 -1737
rect -2248 -1885 -2242 -1833
rect -2190 -1834 -2184 -1833
rect -1610 -1834 -1560 -1780
rect -1306 -1804 -1218 -1777
rect -521 -1727 -8 -1726
rect -521 -1777 -76 -1727
rect -26 -1777 -8 -1727
rect -798 -1834 -792 -1833
rect -2190 -1884 -792 -1834
rect -2190 -1885 -2184 -1884
rect -798 -1885 -792 -1884
rect -740 -1834 -734 -1833
rect -521 -1834 -470 -1777
rect -94 -1796 -8 -1777
rect 493 -1743 551 -1737
rect 917 -1743 951 -1658
rect 1950 -1722 1984 -1658
rect 493 -1777 505 -1743
rect 539 -1777 951 -1743
rect 1456 -1737 1532 -1724
rect 1456 -1777 1479 -1737
rect 1513 -1777 1532 -1737
rect 493 -1783 551 -1777
rect 1456 -1800 1532 -1777
rect 1936 -1737 1996 -1722
rect 2519 -1733 2553 -1612
rect 2892 -1646 2944 -1640
rect 1936 -1777 1950 -1737
rect 1984 -1777 1996 -1737
rect 1936 -1788 1996 -1777
rect 2513 -1736 2559 -1733
rect 2897 -1736 2938 -1646
rect 3300 -1736 3366 -1722
rect 2513 -1737 3366 -1736
rect 2513 -1745 3314 -1737
rect 2513 -1779 2519 -1745
rect 2553 -1777 3314 -1745
rect 3348 -1777 3366 -1737
rect 2553 -1779 2559 -1777
rect 2513 -1791 2559 -1779
rect 3300 -1790 3366 -1777
rect 4082 -1738 4154 -1720
rect 4082 -1778 4102 -1738
rect 4138 -1778 4480 -1738
rect 4082 -1794 4154 -1778
rect -740 -1884 -469 -1834
rect 1479 -1856 1514 -1800
rect 2744 -1856 2750 -1847
rect -740 -1885 -734 -1884
rect 1479 -1891 2750 -1856
rect 1479 -1894 1514 -1891
rect 2744 -1899 2750 -1891
rect 2802 -1899 2808 -1847
rect -3162 -1978 -2343 -1945
rect -931 -1976 -249 -1945
rect 523 -1976 1149 -1945
rect -3162 -2009 -2329 -1978
rect -913 -2007 -259 -1976
rect 549 -1986 1149 -1976
rect 2593 -1986 3248 -1945
rect -897 -2009 -262 -2007
rect 549 -2009 3297 -1986
rect -3162 -2040 -2331 -2009
rect -921 -2040 -185 -2009
rect 534 -2017 3297 -2009
rect 534 -2040 1191 -2017
rect 2593 -2039 3279 -2017
rect -3162 -3042 -3066 -2040
rect -2664 -2256 -2568 -2250
rect -798 -2338 -792 -2286
rect -740 -2338 -734 -2286
rect -2664 -2498 -2568 -2352
rect -2664 -2512 -2487 -2498
rect -2664 -2594 -2461 -2512
rect -1768 -2808 -1694 -2788
rect -2370 -2831 -2282 -2816
rect -2370 -2832 -2352 -2831
rect -2787 -2875 -2352 -2832
rect -2301 -2875 -2282 -2831
rect -1768 -2844 -1748 -2808
rect -1710 -2818 -1694 -2808
rect -1710 -2835 -1440 -2818
rect -1710 -2844 -1511 -2835
rect -1768 -2862 -1511 -2844
rect -2370 -2900 -2282 -2875
rect -1532 -2875 -1511 -2862
rect -1461 -2836 -1440 -2835
rect -791 -2836 -741 -2338
rect -1461 -2875 -741 -2836
rect -1532 -2898 -1440 -2875
rect -3162 -3105 -2458 -3042
rect -3162 -3129 -2459 -3105
rect -3162 -3138 -2475 -3129
<< via1 >>
rect -2664 1088 -2568 1184
rect -2664 490 -2568 586
rect -828 92 -776 144
rect -2664 -358 -2568 -262
rect -828 -246 -776 -194
rect -2242 -478 -2190 -426
rect 2751 -388 2803 -336
rect -1202 -500 -1150 -448
rect -533 -487 -481 -435
rect 2011 -498 2063 -446
rect -1202 -832 -1150 -780
rect 2290 -832 2342 -780
rect -2664 -934 -2568 -838
rect 2893 -1260 2945 -1208
rect -1966 -1344 -1914 -1292
rect -1967 -1632 -1915 -1580
rect -1285 -1598 -1233 -1546
rect -2664 -1826 -2568 -1730
rect 2510 -1612 2562 -1560
rect -2242 -1885 -2190 -1833
rect -792 -1885 -740 -1833
rect 2892 -1640 2944 -1588
rect 2750 -1899 2802 -1847
rect -2664 -2352 -2568 -2256
rect -792 -2338 -740 -2286
<< metal2 >>
rect -2664 1184 -2568 1190
rect -2664 586 -2568 1088
rect -2670 490 -2664 586
rect -2568 490 -2562 586
rect -828 144 -776 150
rect -828 86 -776 92
rect -824 -194 -780 86
rect -834 -246 -828 -194
rect -776 -246 -770 -194
rect -2664 -262 -2568 -256
rect -2664 -838 -2568 -358
rect 2751 -336 2803 -330
rect 2751 -394 2803 -388
rect -2242 -426 -2190 -420
rect -2242 -484 -2190 -478
rect -2670 -934 -2664 -838
rect -2568 -934 -2562 -838
rect -2664 -1730 -2568 -1724
rect -2664 -2256 -2568 -1826
rect -2241 -1827 -2191 -484
rect -1208 -500 -1202 -448
rect -1150 -500 -1144 -448
rect -539 -487 -533 -435
rect -481 -487 -475 -435
rect -1199 -774 -1153 -500
rect -1202 -780 -1150 -774
rect -1202 -838 -1150 -832
rect -1284 -1238 -1233 -1237
rect -532 -1238 -481 -487
rect 2005 -498 2011 -446
rect 2063 -498 2069 -446
rect 2020 -1133 2054 -498
rect 2290 -780 2342 -774
rect 2759 -783 2794 -394
rect 2342 -829 2794 -783
rect 2290 -838 2342 -832
rect 2020 -1167 2553 -1133
rect -1966 -1292 -1914 -1286
rect -1966 -1350 -1914 -1344
rect -1284 -1289 -481 -1238
rect -1961 -1580 -1920 -1350
rect -1284 -1546 -1233 -1289
rect -1973 -1632 -1967 -1580
rect -1915 -1632 -1909 -1580
rect -1291 -1598 -1285 -1546
rect -1233 -1598 -1227 -1546
rect 2519 -1554 2553 -1167
rect 2510 -1560 2562 -1554
rect 2510 -1618 2562 -1612
rect -2242 -1833 -2190 -1827
rect -2242 -1891 -2190 -1885
rect -792 -1833 -740 -1827
rect 2759 -1841 2794 -829
rect 2893 -1208 2945 -1202
rect 2893 -1266 2945 -1260
rect 2898 -1588 2939 -1266
rect 2886 -1640 2892 -1588
rect 2944 -1640 2950 -1588
rect -792 -1891 -740 -1885
rect 2750 -1847 2802 -1841
rect -2670 -2352 -2664 -2256
rect -2568 -2352 -2562 -2256
rect -791 -2280 -741 -1891
rect 2750 -1905 2802 -1899
rect -792 -2286 -740 -2280
rect -792 -2344 -740 -2338
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -2862 0 1 -1992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1704896540
transform 1 0 -2858 0 1 -592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1704896540
transform 1 0 -2664 0 1 -3090
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1704896540
transform 1 0 -2662 0 1 808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_8  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -2494 0 1 808
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x2
timestamp 1704896540
transform 1 0 -2362 0 1 -592
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x3
timestamp 1704896540
transform 1 0 -2362 0 1 -1992
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x4
timestamp 1704896540
transform 1 0 -2504 0 1 -3090
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  x5 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -264 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x6
timestamp 1704896540
transform 1 0 -262 0 1 -1992
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  x7 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1140 0 1 -592
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  x8
timestamp 1704896540
transform 1 0 1138 0 1 -1992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  x9 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3236 0 1 -1992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x10
timestamp 1704896540
transform 1 0 3238 0 1 -592
box -38 -48 1142 592
<< labels >>
rlabel metal1 -2664 -262 -2568 490 7 VPWR
rlabel metal1 -3162 -3138 -3066 856 7 VGND
rlabel metal1 4142 -386 4491 -340 3 Qn
rlabel metal1 4138 -1778 4480 -1738 3 Q
rlabel metal1 -2787 -2875 -2352 -2832 7 ENABLE
rlabel metal1 -2921 922 -2124 972 7 ENABLE
<< end >>
