VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_relax_2
  CLASS BLOCK ;
  FOREIGN tt_um_relax_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT 79.065 105.675 79.395 106.475 ;
        RECT 79.905 105.675 80.235 106.475 ;
        RECT 80.745 105.675 81.075 106.475 ;
        RECT 81.585 105.675 81.915 106.475 ;
        RECT 82.425 105.675 82.755 106.475 ;
        RECT 83.265 105.675 83.595 106.475 ;
        RECT 84.105 105.675 84.435 106.475 ;
        RECT 84.945 105.675 85.275 106.475 ;
        RECT 79.065 105.475 85.275 105.675 ;
        RECT 82.190 105.085 82.670 105.475 ;
        RECT 82.840 105.085 84.855 105.285 ;
        RECT 82.425 104.915 82.670 105.085 ;
        RECT 85.025 104.915 85.275 105.475 ;
        RECT 82.425 104.665 85.275 104.915 ;
        RECT 79.725 98.675 80.055 99.475 ;
        RECT 80.565 98.675 80.895 99.475 ;
        RECT 81.405 98.675 81.735 99.475 ;
        RECT 82.245 98.675 82.575 99.475 ;
        RECT 83.085 98.675 83.415 99.475 ;
        RECT 83.925 98.675 84.255 99.475 ;
        RECT 84.765 98.675 85.095 99.475 ;
        RECT 85.605 98.675 85.935 99.475 ;
        RECT 79.725 98.475 85.935 98.675 ;
        RECT 82.850 98.085 83.330 98.475 ;
        RECT 83.085 97.915 83.330 98.085 ;
        RECT 85.685 97.915 85.935 98.475 ;
        RECT 90.380 98.085 93.235 98.335 ;
        RECT 83.085 97.665 85.935 97.915 ;
        RECT 83.500 91.085 85.515 91.285 ;
      LAYER met1 ;
        RECT 82.220 105.420 82.620 105.580 ;
        RECT 83.030 105.420 83.420 105.470 ;
        RECT 82.220 105.290 83.420 105.420 ;
        RECT 82.220 105.260 87.120 105.290 ;
        RECT 82.220 105.180 82.620 105.260 ;
        RECT 83.030 105.085 87.120 105.260 ;
        RECT 83.030 105.020 83.420 105.085 ;
        RECT 86.900 103.170 87.120 105.085 ;
        RECT 90.370 103.170 91.270 103.200 ;
        RECT 86.900 102.270 91.270 103.170 ;
        RECT 86.900 100.690 87.120 102.270 ;
        RECT 90.370 102.240 91.270 102.270 ;
        RECT 86.850 100.430 87.170 100.690 ;
        RECT 86.880 98.980 87.140 99.030 ;
        RECT 82.950 98.760 88.610 98.980 ;
        RECT 82.950 98.530 83.170 98.760 ;
        RECT 86.880 98.710 87.140 98.760 ;
        RECT 82.830 98.070 83.290 98.530 ;
        RECT 88.355 98.340 88.610 98.760 ;
        RECT 90.500 98.340 90.990 98.460 ;
        RECT 88.355 98.085 90.990 98.340 ;
        RECT 88.355 97.825 88.610 98.085 ;
        RECT 90.500 97.990 90.990 98.085 ;
        RECT 88.355 97.505 88.615 97.825 ;
        RECT 84.595 91.950 84.855 92.270 ;
        RECT 84.595 91.400 84.850 91.950 ;
        RECT 84.490 90.950 84.930 91.400 ;
      LAYER met2 ;
        RECT 99.595 103.170 100.445 103.190 ;
        RECT 90.340 102.270 100.470 103.170 ;
        RECT 99.595 102.250 100.445 102.270 ;
        RECT 86.880 100.400 87.140 100.720 ;
        RECT 86.900 99.000 87.120 100.400 ;
        RECT 86.850 98.740 87.170 99.000 ;
        RECT 88.325 97.535 88.645 97.795 ;
        RECT 84.600 93.780 84.855 93.785 ;
        RECT 88.360 93.780 88.615 97.535 ;
        RECT 84.600 93.525 88.615 93.780 ;
        RECT 84.600 92.240 84.855 93.525 ;
        RECT 84.565 91.980 84.885 92.240 ;
      LAYER met3 ;
        RECT 99.570 102.270 152.710 103.170 ;
        RECT 151.810 4.605 152.710 102.270 ;
        RECT 151.785 3.715 152.735 4.605 ;
        RECT 151.810 3.710 152.710 3.715 ;
      LAYER met4 ;
        RECT 151.810 0.000 152.710 4.610 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT 79.720 98.085 82.575 98.305 ;
        RECT 79.725 91.675 80.055 92.475 ;
        RECT 80.565 91.675 80.895 92.475 ;
        RECT 81.405 91.675 81.735 92.475 ;
        RECT 82.245 91.675 82.575 92.475 ;
        RECT 83.085 91.675 83.415 92.475 ;
        RECT 83.925 91.675 84.255 92.475 ;
        RECT 84.765 91.675 85.095 92.475 ;
        RECT 85.605 91.675 85.935 92.475 ;
        RECT 79.725 91.475 85.935 91.675 ;
        RECT 82.850 91.085 83.330 91.475 ;
        RECT 83.085 90.915 83.330 91.085 ;
        RECT 85.685 90.915 85.935 91.475 ;
        RECT 90.390 91.085 93.245 91.335 ;
        RECT 83.085 90.665 85.935 90.915 ;
        RECT 79.015 86.185 79.345 86.985 ;
        RECT 79.855 86.185 80.185 86.985 ;
        RECT 80.695 86.185 81.025 86.985 ;
        RECT 81.535 86.185 81.865 86.985 ;
        RECT 82.375 86.185 82.705 86.985 ;
        RECT 83.215 86.185 83.545 86.985 ;
        RECT 84.055 86.185 84.385 86.985 ;
        RECT 84.895 86.185 85.225 86.985 ;
        RECT 79.015 85.985 85.225 86.185 ;
        RECT 82.140 85.595 82.620 85.985 ;
        RECT 82.790 85.595 84.805 85.795 ;
        RECT 82.375 85.425 82.620 85.595 ;
        RECT 84.975 85.425 85.225 85.985 ;
        RECT 82.375 85.175 85.225 85.425 ;
      LAYER met1 ;
        RECT 79.815 97.840 80.065 98.335 ;
        RECT 79.780 97.580 80.100 97.840 ;
        RECT 82.850 91.070 83.320 91.520 ;
        RECT 90.550 91.340 90.980 91.420 ;
        RECT 88.415 91.085 90.980 91.340 ;
        RECT 79.780 90.800 80.100 90.805 ;
        RECT 82.970 90.800 83.220 91.070 ;
        RECT 87.030 90.800 87.350 90.805 ;
        RECT 88.415 90.800 88.670 91.085 ;
        RECT 90.550 90.990 90.980 91.085 ;
        RECT 79.780 90.550 88.675 90.800 ;
        RECT 79.780 90.545 80.100 90.550 ;
        RECT 87.030 90.545 87.350 90.550 ;
        RECT 87.030 88.280 87.350 88.540 ;
        RECT 87.065 87.460 87.315 88.280 ;
        RECT 90.010 87.460 90.910 87.490 ;
        RECT 87.065 86.560 90.910 87.460 ;
        RECT 82.180 85.880 82.550 86.030 ;
        RECT 82.180 85.790 83.820 85.880 ;
        RECT 87.065 85.790 87.315 86.560 ;
        RECT 90.010 86.530 90.910 86.560 ;
        RECT 82.180 85.660 87.315 85.790 ;
        RECT 83.360 85.595 87.315 85.660 ;
        RECT 83.360 85.480 83.820 85.595 ;
      LAYER met2 ;
        RECT 79.810 97.550 80.070 97.870 ;
        RECT 79.815 90.835 80.065 97.550 ;
        RECT 79.810 90.515 80.070 90.835 ;
        RECT 87.060 90.515 87.320 90.835 ;
        RECT 87.065 88.570 87.315 90.515 ;
        RECT 87.060 88.250 87.320 88.570 ;
        RECT 89.980 87.435 97.130 87.460 ;
        RECT 89.980 86.585 97.150 87.435 ;
        RECT 89.980 86.560 97.130 86.585 ;
      LAYER met3 ;
        RECT 96.230 86.560 133.390 87.460 ;
        RECT 132.490 5.295 133.390 86.560 ;
        RECT 132.465 4.405 133.415 5.295 ;
        RECT 132.490 4.400 133.390 4.405 ;
      LAYER met4 ;
        RECT 132.490 0.000 133.390 5.300 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 109.055 91.625 109.225 92.475 ;
        RECT 109.895 91.625 110.065 92.475 ;
        RECT 110.735 91.625 110.905 92.475 ;
        RECT 111.575 91.625 111.745 92.475 ;
        RECT 109.055 91.455 111.745 91.625 ;
        RECT 111.490 90.915 111.745 91.455 ;
        RECT 109.055 90.745 111.745 90.915 ;
        RECT 109.055 90.265 109.225 90.745 ;
        RECT 109.895 90.265 110.065 90.745 ;
        RECT 110.735 90.265 110.905 90.745 ;
        RECT 111.575 90.265 111.745 90.745 ;
      LAYER met1 ;
        RECT 116.230 105.610 116.530 105.640 ;
        RECT 115.180 105.310 116.530 105.610 ;
        RECT 111.430 91.280 111.790 91.370 ;
        RECT 115.180 91.280 115.380 105.310 ;
        RECT 116.230 105.280 116.530 105.310 ;
        RECT 111.430 91.080 115.380 91.280 ;
        RECT 111.430 91.000 111.790 91.080 ;
      LAYER met2 ;
        RECT 116.230 113.900 116.530 113.910 ;
        RECT 116.195 113.620 116.565 113.900 ;
        RECT 116.230 105.610 116.530 113.620 ;
        RECT 116.200 105.310 116.560 105.610 ;
      LAYER met3 ;
        RECT 116.190 192.300 116.570 192.620 ;
        RECT 116.230 113.925 116.530 192.300 ;
        RECT 116.215 113.595 116.545 113.925 ;
      LAYER met4 ;
        RECT 116.230 192.625 116.530 225.760 ;
        RECT 116.215 192.295 116.545 192.625 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 109.065 98.625 109.235 99.475 ;
        RECT 109.905 98.625 110.075 99.475 ;
        RECT 110.745 98.625 110.915 99.475 ;
        RECT 111.585 98.625 111.755 99.475 ;
        RECT 109.065 98.455 111.755 98.625 ;
        RECT 111.500 97.915 111.755 98.455 ;
        RECT 109.065 97.745 111.755 97.915 ;
        RECT 109.065 97.265 109.235 97.745 ;
        RECT 109.905 97.265 110.075 97.745 ;
        RECT 110.745 97.265 110.915 97.745 ;
        RECT 111.585 97.265 111.755 97.745 ;
      LAYER met1 ;
        RECT 113.440 105.465 114.065 105.470 ;
        RECT 113.440 105.170 114.295 105.465 ;
        RECT 111.400 98.270 111.830 98.380 ;
        RECT 114.065 98.270 114.295 105.170 ;
        RECT 111.400 98.040 114.295 98.270 ;
        RECT 111.400 97.950 111.830 98.040 ;
      LAYER met2 ;
        RECT 113.470 113.860 113.770 113.870 ;
        RECT 113.435 113.580 113.805 113.860 ;
        RECT 113.470 105.140 113.770 113.580 ;
      LAYER met3 ;
        RECT 113.460 190.430 113.780 190.810 ;
        RECT 113.470 113.885 113.770 190.430 ;
        RECT 113.455 113.555 113.785 113.885 ;
      LAYER met4 ;
        RECT 113.470 190.785 113.770 225.760 ;
        RECT 113.455 190.455 113.785 190.785 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 79.060 105.085 81.915 105.305 ;
      LAYER met1 ;
        RECT 76.665 108.245 80.630 108.250 ;
        RECT 76.415 107.950 80.630 108.245 ;
        RECT 76.415 104.830 76.665 107.950 ;
        RECT 80.050 104.990 80.480 105.380 ;
        RECT 80.150 104.830 80.400 104.990 ;
        RECT 76.415 104.580 80.400 104.830 ;
      LAYER met2 ;
        RECT 80.310 110.560 80.590 110.595 ;
        RECT 80.300 107.920 80.600 110.560 ;
      LAYER met3 ;
        RECT 110.700 190.500 111.020 190.540 ;
        RECT 80.300 190.200 111.020 190.500 ;
        RECT 80.300 110.575 80.600 190.200 ;
        RECT 110.700 190.160 111.020 190.200 ;
        RECT 80.285 110.245 80.615 110.575 ;
      LAYER met4 ;
        RECT 110.710 190.515 111.010 225.760 ;
        RECT 110.695 190.185 111.025 190.515 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 79.010 85.595 81.865 85.815 ;
      LAYER met1 ;
        RECT 76.635 85.810 76.955 85.835 ;
        RECT 79.170 85.810 79.610 85.890 ;
        RECT 76.635 85.595 79.610 85.810 ;
        RECT 76.635 85.575 76.955 85.595 ;
        RECT 79.170 85.470 79.610 85.595 ;
      LAYER met2 ;
        RECT 74.800 127.950 75.100 127.960 ;
        RECT 74.765 127.670 75.135 127.950 ;
        RECT 73.105 112.280 73.320 112.285 ;
        RECT 74.800 112.280 75.100 127.670 ;
        RECT 73.105 111.980 75.100 112.280 ;
        RECT 73.105 85.815 73.320 111.980 ;
        RECT 76.665 85.815 76.925 85.865 ;
        RECT 73.105 85.600 76.925 85.815 ;
        RECT 76.665 85.545 76.925 85.600 ;
      LAYER met3 ;
        RECT 107.940 197.580 108.260 197.620 ;
        RECT 74.800 197.280 108.260 197.580 ;
        RECT 74.800 127.975 75.100 197.280 ;
        RECT 107.940 197.240 108.260 197.280 ;
        RECT 74.785 127.645 75.115 127.975 ;
      LAYER met4 ;
        RECT 107.950 197.595 108.250 225.760 ;
        RECT 107.935 197.265 108.265 197.595 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 77.520 105.315 86.100 106.920 ;
        RECT 76.540 98.315 112.920 99.920 ;
        RECT 76.520 91.315 112.910 92.920 ;
        RECT 106.130 91.305 106.970 91.315 ;
        RECT 77.090 87.420 86.050 87.430 ;
        RECT 76.860 85.825 86.050 87.420 ;
        RECT 76.860 85.815 77.700 85.825 ;
      LAYER li1 ;
        RECT 77.710 106.645 78.170 106.815 ;
        RECT 78.550 106.645 85.910 106.815 ;
        RECT 77.795 105.480 78.085 106.645 ;
        RECT 78.640 105.505 78.895 106.645 ;
        RECT 79.565 105.845 79.735 106.645 ;
        RECT 80.405 105.845 80.575 106.645 ;
        RECT 81.245 105.845 81.415 106.645 ;
        RECT 82.085 105.845 82.255 106.645 ;
        RECT 82.925 105.845 83.095 106.645 ;
        RECT 83.765 105.845 83.935 106.645 ;
        RECT 84.605 105.845 84.775 106.645 ;
        RECT 85.465 105.505 85.820 106.645 ;
        RECT 76.730 99.645 77.190 99.815 ;
        RECT 79.210 99.645 86.570 99.815 ;
        RECT 89.700 99.645 93.840 99.815 ;
        RECT 96.720 99.645 104.080 99.815 ;
        RECT 105.660 99.645 106.120 99.815 ;
        RECT 107.210 99.645 112.730 99.815 ;
        RECT 76.815 98.480 77.105 99.645 ;
        RECT 79.300 98.505 79.555 99.645 ;
        RECT 80.225 98.845 80.395 99.645 ;
        RECT 81.065 98.845 81.235 99.645 ;
        RECT 81.905 98.845 82.075 99.645 ;
        RECT 82.745 98.845 82.915 99.645 ;
        RECT 83.585 98.845 83.755 99.645 ;
        RECT 84.425 98.845 84.595 99.645 ;
        RECT 85.265 98.845 85.435 99.645 ;
        RECT 86.125 98.505 86.480 99.645 ;
        RECT 89.955 98.845 90.210 99.645 ;
        RECT 90.880 98.845 91.050 99.645 ;
        RECT 91.720 98.845 91.890 99.645 ;
        RECT 92.560 98.845 92.730 99.645 ;
        RECT 93.400 98.845 93.700 99.645 ;
        RECT 97.295 98.845 97.545 99.645 ;
        RECT 98.135 98.845 98.385 99.645 ;
        RECT 98.975 98.845 99.225 99.645 ;
        RECT 99.815 98.845 100.065 99.645 ;
        RECT 105.745 98.480 106.035 99.645 ;
        RECT 107.805 98.845 107.975 99.645 ;
        RECT 108.645 98.845 108.815 99.645 ;
        RECT 109.405 98.845 109.735 99.645 ;
        RECT 110.245 98.845 110.575 99.645 ;
        RECT 111.085 98.845 111.415 99.645 ;
        RECT 111.925 98.495 112.255 99.645 ;
        RECT 76.710 92.645 77.170 92.815 ;
        RECT 79.210 92.645 86.570 92.815 ;
        RECT 89.710 92.645 93.850 92.815 ;
        RECT 96.710 92.645 104.070 92.815 ;
        RECT 76.795 91.480 77.085 92.645 ;
        RECT 79.300 91.505 79.555 92.645 ;
        RECT 80.225 91.845 80.395 92.645 ;
        RECT 81.065 91.845 81.235 92.645 ;
        RECT 81.905 91.845 82.075 92.645 ;
        RECT 82.745 91.845 82.915 92.645 ;
        RECT 83.585 91.845 83.755 92.645 ;
        RECT 84.425 91.845 84.595 92.645 ;
        RECT 85.265 91.845 85.435 92.645 ;
        RECT 86.125 91.505 86.480 92.645 ;
        RECT 89.965 91.845 90.220 92.645 ;
        RECT 90.890 91.845 91.060 92.645 ;
        RECT 91.730 91.845 91.900 92.645 ;
        RECT 92.570 91.845 92.740 92.645 ;
        RECT 93.410 91.845 93.710 92.645 ;
        RECT 97.285 91.845 97.535 92.645 ;
        RECT 98.125 91.845 98.375 92.645 ;
        RECT 98.965 91.845 99.215 92.645 ;
        RECT 99.805 91.845 100.055 92.645 ;
        RECT 106.320 92.635 106.780 92.805 ;
        RECT 107.200 92.645 112.720 92.815 ;
        RECT 106.405 91.470 106.695 92.635 ;
        RECT 107.795 91.845 107.965 92.645 ;
        RECT 108.635 91.845 108.805 92.645 ;
        RECT 109.395 91.845 109.725 92.645 ;
        RECT 110.235 91.845 110.565 92.645 ;
        RECT 111.075 91.845 111.405 92.645 ;
        RECT 111.915 91.495 112.245 92.645 ;
        RECT 77.050 87.145 77.510 87.315 ;
        RECT 78.500 87.155 85.860 87.325 ;
        RECT 77.135 85.980 77.425 87.145 ;
        RECT 78.590 86.015 78.845 87.155 ;
        RECT 79.515 86.355 79.685 87.155 ;
        RECT 80.355 86.355 80.525 87.155 ;
        RECT 81.195 86.355 81.365 87.155 ;
        RECT 82.035 86.355 82.205 87.155 ;
        RECT 82.875 86.355 83.045 87.155 ;
        RECT 83.715 86.355 83.885 87.155 ;
        RECT 84.555 86.355 84.725 87.155 ;
        RECT 85.415 86.015 85.770 87.155 ;
      LAYER met1 ;
        RECT 77.710 106.870 85.910 106.970 ;
        RECT 77.700 106.490 85.910 106.870 ;
        RECT 77.700 105.890 78.180 106.490 ;
        RECT 77.670 105.410 78.210 105.890 ;
        RECT 77.700 102.240 78.180 102.930 ;
        RECT 76.490 101.760 78.180 102.240 ;
        RECT 77.700 99.970 78.180 101.760 ;
        RECT 76.730 99.490 112.730 99.970 ;
        RECT 77.700 98.660 78.180 99.490 ;
        RECT 77.670 98.180 78.210 98.660 ;
        RECT 77.700 92.970 78.180 95.810 ;
        RECT 76.710 92.495 112.720 92.970 ;
        RECT 76.710 92.490 77.170 92.495 ;
        RECT 77.700 91.320 78.180 92.495 ;
        RECT 79.210 92.490 86.570 92.495 ;
        RECT 89.710 92.490 93.850 92.495 ;
        RECT 96.710 92.490 104.070 92.495 ;
        RECT 106.320 92.480 106.780 92.495 ;
        RECT 107.200 92.490 112.720 92.495 ;
        RECT 77.670 90.840 78.210 91.320 ;
        RECT 77.670 88.310 78.210 88.790 ;
        RECT 77.700 87.470 78.180 88.310 ;
        RECT 78.500 87.470 85.860 87.480 ;
        RECT 77.050 87.000 85.860 87.470 ;
        RECT 77.050 86.990 77.510 87.000 ;
      LAYER met2 ;
        RECT 77.700 102.900 78.180 105.920 ;
        RECT 77.670 102.420 78.210 102.900 ;
        RECT 76.520 102.240 77.000 102.270 ;
        RECT 73.885 101.760 77.000 102.240 ;
        RECT 76.520 101.730 77.000 101.760 ;
        RECT 77.700 95.780 78.180 98.690 ;
        RECT 77.670 95.300 78.210 95.780 ;
        RECT 77.700 88.280 78.180 91.350 ;
      LAYER met3 ;
        RECT 73.905 102.240 74.435 102.265 ;
        RECT 69.350 101.760 74.435 102.240 ;
        RECT 1.000 100.430 31.105 100.710 ;
        RECT 69.385 100.430 70.795 101.760 ;
        RECT 73.905 101.735 74.435 101.760 ;
        RECT 1.000 99.020 70.795 100.430 ;
        RECT 1.000 98.740 31.105 99.020 ;
        RECT 1.000 98.710 3.000 98.740 ;
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 77.715 104.115 85.905 105.025 ;
        RECT 78.700 103.925 78.870 104.115 ;
        RECT 76.725 97.115 112.345 98.025 ;
        RECT 79.360 96.925 79.530 97.115 ;
        RECT 89.870 97.095 90.015 97.115 ;
        RECT 89.845 96.925 90.015 97.095 ;
        RECT 96.865 96.925 97.035 97.115 ;
        RECT 107.360 96.925 107.530 97.115 ;
        RECT 76.725 90.115 112.335 91.025 ;
        RECT 79.360 89.925 79.530 90.115 ;
        RECT 89.880 90.095 90.025 90.115 ;
        RECT 89.855 89.925 90.025 90.095 ;
        RECT 96.855 89.925 97.025 90.115 ;
        RECT 107.350 89.925 107.520 90.115 ;
        RECT 77.045 84.625 85.855 85.535 ;
        RECT 78.650 84.435 78.820 84.625 ;
      LAYER li1 ;
        RECT 77.795 104.095 78.085 104.820 ;
        RECT 79.145 104.095 79.315 104.575 ;
        RECT 79.985 104.095 80.155 104.575 ;
        RECT 80.825 104.095 80.995 104.575 ;
        RECT 81.665 104.095 81.835 104.575 ;
        RECT 77.710 103.925 78.170 104.095 ;
        RECT 78.550 103.925 85.910 104.095 ;
        RECT 76.815 97.095 77.105 97.820 ;
        RECT 79.805 97.095 79.975 97.575 ;
        RECT 80.645 97.095 80.815 97.575 ;
        RECT 81.485 97.095 81.655 97.575 ;
        RECT 82.325 97.095 82.495 97.575 ;
        RECT 89.955 97.095 90.210 97.555 ;
        RECT 90.880 97.095 91.050 97.555 ;
        RECT 91.720 97.095 91.890 97.555 ;
        RECT 92.560 97.095 92.730 97.555 ;
        RECT 93.400 97.095 93.705 97.555 ;
        RECT 96.810 97.095 97.085 97.915 ;
        RECT 97.755 97.095 97.925 97.565 ;
        RECT 98.595 97.095 98.765 97.565 ;
        RECT 99.435 97.095 99.605 97.565 ;
        RECT 100.275 97.095 100.445 97.565 ;
        RECT 101.115 97.095 101.285 97.565 ;
        RECT 101.955 97.095 102.125 97.565 ;
        RECT 102.795 97.095 102.965 97.565 ;
        RECT 103.635 97.095 103.925 97.565 ;
        RECT 105.745 97.095 106.035 97.820 ;
        RECT 107.725 97.095 108.055 97.575 ;
        RECT 108.565 97.095 108.895 97.575 ;
        RECT 109.405 97.095 109.735 97.575 ;
        RECT 110.245 97.095 110.575 97.575 ;
        RECT 111.085 97.095 111.415 97.575 ;
        RECT 111.925 97.095 112.255 97.895 ;
        RECT 76.730 96.925 77.190 97.095 ;
        RECT 79.210 96.925 86.570 97.095 ;
        RECT 89.700 96.925 93.840 97.095 ;
        RECT 96.720 96.925 104.080 97.095 ;
        RECT 105.660 96.925 106.120 97.095 ;
        RECT 107.210 96.925 112.730 97.095 ;
        RECT 76.795 90.095 77.085 90.820 ;
        RECT 79.805 90.095 79.975 90.575 ;
        RECT 80.645 90.095 80.815 90.575 ;
        RECT 81.485 90.095 81.655 90.575 ;
        RECT 82.325 90.095 82.495 90.575 ;
        RECT 89.965 90.095 90.220 90.555 ;
        RECT 90.890 90.095 91.060 90.555 ;
        RECT 91.730 90.095 91.900 90.555 ;
        RECT 92.570 90.095 92.740 90.555 ;
        RECT 93.410 90.095 93.715 90.555 ;
        RECT 96.800 90.095 97.075 90.915 ;
        RECT 97.745 90.095 97.915 90.565 ;
        RECT 98.585 90.095 98.755 90.565 ;
        RECT 99.425 90.095 99.595 90.565 ;
        RECT 100.265 90.095 100.435 90.565 ;
        RECT 101.105 90.095 101.275 90.565 ;
        RECT 101.945 90.095 102.115 90.565 ;
        RECT 102.785 90.095 102.955 90.565 ;
        RECT 103.625 90.095 103.915 90.565 ;
        RECT 76.710 89.925 77.170 90.095 ;
        RECT 79.210 89.925 86.570 90.095 ;
        RECT 89.710 89.925 93.850 90.095 ;
        RECT 96.710 89.925 104.070 90.095 ;
        RECT 106.405 90.085 106.695 90.810 ;
        RECT 107.715 90.095 108.045 90.575 ;
        RECT 108.555 90.095 108.885 90.575 ;
        RECT 109.395 90.095 109.725 90.575 ;
        RECT 110.235 90.095 110.565 90.575 ;
        RECT 111.075 90.095 111.405 90.575 ;
        RECT 111.915 90.095 112.245 90.895 ;
        RECT 106.320 89.915 106.780 90.085 ;
        RECT 107.200 89.925 112.720 90.095 ;
        RECT 77.135 84.595 77.425 85.320 ;
        RECT 79.095 84.605 79.265 85.085 ;
        RECT 79.935 84.605 80.105 85.085 ;
        RECT 80.775 84.605 80.945 85.085 ;
        RECT 81.615 84.605 81.785 85.085 ;
        RECT 77.050 84.425 77.510 84.595 ;
        RECT 78.500 84.435 85.860 84.605 ;
      LAYER met1 ;
        RECT 72.480 103.770 85.910 104.250 ;
        RECT 72.480 97.250 72.960 103.770 ;
        RECT 72.480 96.770 112.730 97.250 ;
        RECT 72.480 90.245 72.960 96.770 ;
        RECT 76.710 90.245 77.170 90.250 ;
        RECT 79.210 90.245 86.570 90.250 ;
        RECT 89.710 90.245 93.850 90.250 ;
        RECT 96.710 90.245 104.070 90.250 ;
        RECT 107.200 90.245 112.720 90.250 ;
        RECT 58.710 90.210 60.710 90.240 ;
        RECT 72.480 90.210 112.720 90.245 ;
        RECT 58.710 89.775 112.720 90.210 ;
        RECT 58.710 89.770 104.070 89.775 ;
        RECT 58.710 88.210 72.960 89.770 ;
        RECT 106.320 89.760 106.780 89.775 ;
        RECT 107.200 89.770 112.720 89.775 ;
        RECT 58.710 88.180 60.710 88.210 ;
        RECT 72.480 84.760 72.960 88.210 ;
        RECT 72.480 84.280 85.860 84.760 ;
        RECT 72.480 84.260 72.960 84.280 ;
        RECT 77.050 84.270 77.510 84.280 ;
      LAYER met2 ;
        RECT 45.025 90.210 46.975 90.230 ;
        RECT 45.000 88.210 60.740 90.210 ;
        RECT 45.025 88.190 46.975 88.210 ;
      LAYER met3 ;
        RECT 15.495 90.210 17.485 90.235 ;
        RECT 15.490 88.210 47.000 90.210 ;
        RECT 15.495 88.185 17.485 88.210 ;
      LAYER met4 ;
        RECT 4.000 90.210 6.000 220.760 ;
        RECT 4.000 88.210 17.490 90.210 ;
        RECT 4.000 5.000 6.000 88.210 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 78.640 104.745 82.255 104.915 ;
        RECT 78.640 104.265 78.975 104.745 ;
        RECT 79.485 104.265 79.815 104.745 ;
        RECT 80.325 104.265 80.655 104.745 ;
        RECT 81.165 104.265 81.495 104.745 ;
        RECT 82.005 104.495 82.255 104.745 ;
        RECT 85.445 104.495 85.820 104.915 ;
        RECT 82.005 104.265 85.820 104.495 ;
        RECT 90.380 98.675 90.710 99.475 ;
        RECT 91.220 98.675 91.550 99.475 ;
        RECT 92.060 98.675 92.390 99.475 ;
        RECT 92.900 98.675 93.230 99.475 ;
        RECT 96.810 98.675 97.125 99.475 ;
        RECT 97.715 98.675 97.965 99.475 ;
        RECT 98.555 98.675 98.805 99.475 ;
        RECT 99.395 98.675 99.645 99.475 ;
        RECT 100.235 99.305 103.845 99.475 ;
        RECT 100.235 98.675 100.485 99.305 ;
        RECT 89.785 98.505 93.755 98.675 ;
        RECT 83.500 98.085 85.515 98.285 ;
        RECT 89.785 97.915 90.130 98.505 ;
        RECT 93.435 97.915 93.755 98.505 ;
        RECT 96.810 98.465 100.485 98.675 ;
        RECT 100.655 98.625 100.905 99.135 ;
        RECT 101.075 98.795 101.325 99.305 ;
        RECT 101.495 98.625 101.745 99.135 ;
        RECT 101.915 98.795 102.165 99.305 ;
        RECT 102.335 98.625 102.585 99.135 ;
        RECT 102.755 98.795 103.005 99.305 ;
        RECT 103.175 98.625 103.425 99.135 ;
        RECT 103.595 98.795 103.845 99.305 ;
        RECT 107.305 98.625 107.635 99.475 ;
        RECT 108.145 98.625 108.475 99.475 ;
        RECT 100.655 98.455 103.995 98.625 ;
        RECT 107.305 98.455 108.805 98.625 ;
        RECT 97.080 98.085 100.250 98.285 ;
        RECT 100.520 98.085 103.260 98.285 ;
        RECT 103.430 97.915 103.995 98.455 ;
        RECT 107.350 98.085 108.450 98.285 ;
        RECT 108.630 98.255 108.805 98.455 ;
        RECT 108.630 98.085 111.255 98.255 ;
        RECT 108.630 97.915 108.805 98.085 ;
        RECT 79.300 97.745 82.915 97.915 ;
        RECT 79.300 97.265 79.635 97.745 ;
        RECT 80.145 97.265 80.475 97.745 ;
        RECT 80.985 97.265 81.315 97.745 ;
        RECT 81.825 97.265 82.155 97.745 ;
        RECT 82.665 97.495 82.915 97.745 ;
        RECT 86.105 97.495 86.480 97.915 ;
        RECT 89.785 97.725 93.755 97.915 ;
        RECT 97.255 97.735 103.995 97.915 ;
        RECT 107.385 97.745 108.805 97.915 ;
        RECT 82.665 97.265 86.480 97.495 ;
        RECT 90.380 97.265 90.710 97.725 ;
        RECT 91.220 97.265 91.550 97.725 ;
        RECT 92.060 97.265 92.390 97.725 ;
        RECT 92.900 97.265 93.230 97.725 ;
        RECT 97.255 97.265 97.585 97.735 ;
        RECT 98.095 97.265 98.425 97.735 ;
        RECT 98.935 97.265 99.265 97.735 ;
        RECT 99.775 97.265 100.105 97.735 ;
        RECT 100.615 97.265 100.945 97.735 ;
        RECT 101.455 97.265 101.785 97.735 ;
        RECT 102.295 97.265 102.625 97.735 ;
        RECT 103.135 97.265 103.465 97.735 ;
        RECT 107.385 97.265 107.555 97.745 ;
        RECT 108.225 97.270 108.395 97.745 ;
        RECT 90.390 91.675 90.720 92.475 ;
        RECT 91.230 91.675 91.560 92.475 ;
        RECT 92.070 91.675 92.400 92.475 ;
        RECT 92.910 91.675 93.240 92.475 ;
        RECT 96.800 91.675 97.115 92.475 ;
        RECT 97.705 91.675 97.955 92.475 ;
        RECT 98.545 91.675 98.795 92.475 ;
        RECT 99.385 91.675 99.635 92.475 ;
        RECT 100.225 92.305 103.835 92.475 ;
        RECT 100.225 91.675 100.475 92.305 ;
        RECT 89.795 91.505 93.765 91.675 ;
        RECT 79.720 91.085 82.575 91.305 ;
        RECT 89.795 90.915 90.140 91.505 ;
        RECT 93.445 90.915 93.765 91.505 ;
        RECT 96.800 91.465 100.475 91.675 ;
        RECT 100.645 91.625 100.895 92.135 ;
        RECT 101.065 91.795 101.315 92.305 ;
        RECT 101.485 91.625 101.735 92.135 ;
        RECT 101.905 91.795 102.155 92.305 ;
        RECT 102.325 91.625 102.575 92.135 ;
        RECT 102.745 91.795 102.995 92.305 ;
        RECT 103.165 91.625 103.415 92.135 ;
        RECT 103.585 91.795 103.835 92.305 ;
        RECT 107.295 91.625 107.625 92.475 ;
        RECT 108.135 91.625 108.465 92.475 ;
        RECT 100.645 91.455 103.985 91.625 ;
        RECT 107.295 91.455 108.795 91.625 ;
        RECT 97.070 91.085 100.240 91.285 ;
        RECT 100.510 91.085 103.250 91.285 ;
        RECT 103.420 90.915 103.985 91.455 ;
        RECT 107.340 91.085 108.440 91.285 ;
        RECT 108.620 91.255 108.795 91.455 ;
        RECT 108.620 91.085 111.245 91.255 ;
        RECT 108.620 90.915 108.795 91.085 ;
        RECT 79.300 90.745 82.915 90.915 ;
        RECT 79.300 90.265 79.635 90.745 ;
        RECT 80.145 90.265 80.475 90.745 ;
        RECT 80.985 90.265 81.315 90.745 ;
        RECT 81.825 90.265 82.155 90.745 ;
        RECT 82.665 90.495 82.915 90.745 ;
        RECT 86.105 90.495 86.480 90.915 ;
        RECT 89.795 90.725 93.765 90.915 ;
        RECT 97.245 90.735 103.985 90.915 ;
        RECT 107.375 90.745 108.795 90.915 ;
        RECT 82.665 90.265 86.480 90.495 ;
        RECT 90.390 90.265 90.720 90.725 ;
        RECT 91.230 90.265 91.560 90.725 ;
        RECT 92.070 90.265 92.400 90.725 ;
        RECT 92.910 90.265 93.240 90.725 ;
        RECT 97.245 90.265 97.575 90.735 ;
        RECT 98.085 90.265 98.415 90.735 ;
        RECT 98.925 90.265 99.255 90.735 ;
        RECT 99.765 90.265 100.095 90.735 ;
        RECT 100.605 90.265 100.935 90.735 ;
        RECT 101.445 90.265 101.775 90.735 ;
        RECT 102.285 90.265 102.615 90.735 ;
        RECT 103.125 90.265 103.455 90.735 ;
        RECT 107.375 90.265 107.545 90.745 ;
        RECT 108.215 90.270 108.385 90.745 ;
        RECT 78.590 85.255 82.205 85.425 ;
        RECT 78.590 84.775 78.925 85.255 ;
        RECT 79.435 84.775 79.765 85.255 ;
        RECT 80.275 84.775 80.605 85.255 ;
        RECT 81.115 84.775 81.445 85.255 ;
        RECT 81.955 85.005 82.205 85.255 ;
        RECT 85.395 85.005 85.770 85.425 ;
        RECT 81.955 84.775 85.770 85.005 ;
      LAYER met1 ;
        RECT 84.920 97.970 85.370 98.390 ;
        RECT 93.450 98.290 93.740 98.305 ;
        RECT 97.630 98.290 98.050 98.350 ;
        RECT 93.450 98.085 98.050 98.290 ;
        RECT 93.450 98.075 93.740 98.085 ;
        RECT 97.630 98.020 98.050 98.085 ;
        RECT 101.030 97.970 101.370 98.350 ;
        RECT 103.640 98.250 103.930 98.280 ;
        RECT 104.745 98.250 105.065 98.290 ;
        RECT 107.510 98.250 107.850 98.370 ;
        RECT 103.640 98.075 107.850 98.250 ;
        RECT 103.640 98.050 103.930 98.075 ;
        RECT 104.745 98.030 105.065 98.075 ;
        RECT 107.510 97.970 107.850 98.075 ;
        RECT 85.025 97.760 85.255 97.970 ;
        RECT 101.120 97.770 101.290 97.970 ;
        RECT 85.010 97.440 85.270 97.760 ;
        RECT 101.075 97.450 101.335 97.770 ;
        RECT 84.980 96.055 85.300 96.070 ;
        RECT 102.440 96.055 102.760 96.070 ;
        RECT 84.980 95.825 102.760 96.055 ;
        RECT 84.980 95.810 85.300 95.825 ;
        RECT 102.440 95.810 102.760 95.825 ;
        RECT 105.455 93.905 105.775 93.930 ;
        RECT 81.220 93.700 105.775 93.905 ;
        RECT 81.220 93.510 81.425 93.700 ;
        RECT 105.455 93.670 105.775 93.700 ;
        RECT 81.160 93.250 81.480 93.510 ;
        RECT 81.185 91.780 81.445 92.100 ;
        RECT 103.540 91.910 103.860 92.170 ;
        RECT 81.210 91.370 81.415 91.780 ;
        RECT 95.605 91.680 100.940 91.850 ;
        RECT 81.140 91.040 81.450 91.370 ;
        RECT 93.485 91.255 93.775 91.285 ;
        RECT 95.605 91.255 95.775 91.680 ;
        RECT 100.770 91.360 100.940 91.680 ;
        RECT 93.485 91.085 95.775 91.255 ;
        RECT 93.485 91.055 93.775 91.085 ;
        RECT 98.300 90.970 98.680 91.350 ;
        RECT 100.700 91.030 101.000 91.360 ;
        RECT 103.615 91.305 103.785 91.910 ;
        RECT 105.480 91.740 105.740 92.060 ;
        RECT 103.585 91.290 103.815 91.305 ;
        RECT 105.505 91.290 105.710 91.740 ;
        RECT 107.520 91.290 107.850 91.360 ;
        RECT 103.585 91.085 107.850 91.290 ;
        RECT 103.585 91.015 103.815 91.085 ;
        RECT 107.520 91.020 107.850 91.085 ;
        RECT 98.415 90.690 98.590 90.970 ;
        RECT 104.740 90.690 105.060 90.735 ;
        RECT 98.415 90.515 105.060 90.690 ;
        RECT 98.415 90.500 98.590 90.515 ;
        RECT 104.740 90.475 105.060 90.515 ;
      LAYER met2 ;
        RECT 104.775 98.000 105.035 98.320 ;
        RECT 84.980 97.470 85.300 97.730 ;
        RECT 101.045 97.480 101.365 97.740 ;
        RECT 85.025 96.100 85.255 97.470 ;
        RECT 85.010 95.780 85.270 96.100 ;
        RECT 101.120 94.305 101.290 97.480 ;
        RECT 102.470 96.055 102.730 96.100 ;
        RECT 104.815 96.055 104.990 98.000 ;
        RECT 102.470 95.825 104.990 96.055 ;
        RECT 102.470 95.780 102.730 95.825 ;
        RECT 101.120 94.135 103.785 94.305 ;
        RECT 81.190 93.220 81.450 93.540 ;
        RECT 81.215 92.070 81.420 93.220 ;
        RECT 103.615 92.200 103.785 94.135 ;
        RECT 81.155 91.810 81.475 92.070 ;
        RECT 103.570 91.880 103.830 92.200 ;
        RECT 104.815 90.765 104.990 95.825 ;
        RECT 105.485 93.640 105.745 93.960 ;
        RECT 105.510 92.030 105.715 93.640 ;
        RECT 105.450 91.770 105.770 92.030 ;
        RECT 104.770 90.445 105.030 90.765 ;
  END
END tt_um_relax_2
END LIBRARY

