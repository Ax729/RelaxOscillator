magic
tech sky130A
magscale 1 2
timestamp 1762226273
<< metal1 >>
rect 15333 21649 16060 21650
rect 15283 21590 16060 21649
rect 16120 21590 16126 21650
rect 15283 20916 15333 21590
rect 23246 21122 23306 21128
rect 22688 21034 22694 21094
rect 22754 21093 22813 21094
rect 22754 21034 22859 21093
rect 18074 20634 18254 20640
rect 17382 20454 18074 20634
rect 18074 20448 18254 20454
rect 15298 20352 15304 20448
rect 15400 20352 15636 20448
rect 22813 19654 22859 21034
rect 22633 19608 22859 19654
rect 23036 21062 23246 21122
rect 23036 18256 23076 21062
rect 23246 21056 23306 21062
rect 22630 18216 23076 18256
rect 11742 18042 12142 18048
rect 12142 17642 14546 18042
rect 11742 17636 12142 17642
rect 15411 17400 15821 17494
rect 18002 17492 18182 17498
rect 17444 17312 18002 17492
rect 18002 17306 18182 17312
rect 15327 17115 15333 17167
rect 15385 17162 15391 17167
rect 15385 17119 15478 17162
rect 15385 17115 15391 17119
<< via1 >>
rect 16060 21590 16120 21650
rect 22694 21034 22754 21094
rect 18074 20454 18254 20634
rect 15304 20352 15400 20448
rect 23246 21062 23306 21122
rect 11742 17642 12142 18042
rect 18002 17312 18182 17492
rect 15333 17115 15385 17167
<< metal2 >>
rect 14960 25590 15020 25592
rect 14953 25534 14962 25590
rect 15018 25534 15027 25590
rect 14621 22456 14664 22457
rect 14960 22456 15020 25534
rect 23246 22780 23306 22782
rect 22694 22772 22754 22774
rect 22687 22716 22696 22772
rect 22752 22716 22761 22772
rect 23239 22724 23248 22780
rect 23304 22724 23313 22780
rect 14621 22396 15020 22456
rect 9005 18042 9395 18046
rect 9000 18037 11742 18042
rect 9000 17647 9005 18037
rect 9395 17647 11742 18037
rect 9000 17642 11742 17647
rect 12142 17642 12148 18042
rect 9005 17638 9395 17642
rect 14621 17163 14664 22396
rect 16062 22112 16118 22119
rect 16060 22110 16120 22112
rect 16060 22054 16062 22110
rect 16118 22054 16120 22110
rect 16060 21650 16120 22054
rect 16060 21584 16120 21590
rect 22694 21094 22754 22716
rect 23246 21122 23306 22724
rect 23240 21062 23246 21122
rect 23306 21062 23312 21122
rect 22694 21028 22754 21034
rect 19919 20634 20089 20638
rect 18068 20454 18074 20634
rect 18254 20629 20094 20634
rect 18254 20459 19919 20629
rect 20089 20459 20094 20629
rect 18254 20454 20094 20459
rect 15304 20448 15400 20454
rect 19919 20450 20089 20454
rect 14777 20352 14786 20448
rect 14882 20352 15304 20448
rect 15304 20346 15400 20352
rect 17996 17312 18002 17492
rect 18182 17487 19426 17492
rect 18182 17317 19251 17487
rect 19421 17317 19430 17487
rect 18182 17312 19426 17317
rect 15333 17167 15385 17173
rect 14621 17120 15333 17163
rect 15333 17109 15385 17115
<< via2 >>
rect 14962 25534 15018 25590
rect 22696 22716 22752 22772
rect 23248 22724 23304 22780
rect 9005 17647 9395 18037
rect 16062 22054 16118 22110
rect 19919 20459 20089 20629
rect 14786 20352 14882 20448
rect 19251 17317 19421 17487
<< metal3 >>
rect 21588 39518 21652 39524
rect 14960 39456 21588 39516
rect 14960 25595 15020 39456
rect 21588 39448 21652 39454
rect 23238 38460 23244 38524
rect 23308 38460 23314 38524
rect 22692 38156 22756 38162
rect 22140 38102 22204 38108
rect 16060 38040 22140 38100
rect 14957 25590 15023 25595
rect 14957 25534 14962 25590
rect 15018 25534 15023 25590
rect 14957 25529 15023 25534
rect 16060 22115 16120 38040
rect 22692 38086 22756 38092
rect 22140 38032 22204 38038
rect 22694 22777 22754 38086
rect 23246 22785 23306 38460
rect 23243 22780 23309 22785
rect 22691 22772 22757 22777
rect 22691 22716 22696 22772
rect 22752 22716 22757 22772
rect 23243 22724 23248 22780
rect 23304 22724 23309 22780
rect 23243 22719 23309 22724
rect 22691 22711 22757 22716
rect 16057 22110 16123 22115
rect 16057 22054 16062 22110
rect 16118 22054 16123 22110
rect 16057 22049 16123 22054
rect 19914 20629 30542 20634
rect 19914 20459 19919 20629
rect 20089 20459 30542 20629
rect 19914 20454 30542 20459
rect 14781 20448 14887 20453
rect 13870 20352 14786 20448
rect 14882 20352 14887 20448
rect 200 20124 6221 20142
rect 200 19758 220 20124
rect 574 20086 6221 20124
rect 13877 20086 14159 20352
rect 14781 20347 14887 20352
rect 574 19804 14159 20086
rect 574 19758 6221 19804
rect 200 19748 6221 19758
rect 200 19742 600 19748
rect 3099 18042 3497 18047
rect 3098 18041 9400 18042
rect 3098 17643 3099 18041
rect 3497 18037 9400 18041
rect 3497 17647 9005 18037
rect 9395 17647 9400 18037
rect 3497 17643 9400 17647
rect 3098 17642 9400 17643
rect 3099 17637 3497 17642
rect 19246 17487 26678 17492
rect 19246 17317 19251 17487
rect 19421 17317 26678 17487
rect 19246 17312 26678 17317
rect 26498 1059 26678 17312
rect 26493 881 26499 1059
rect 26677 881 26683 1059
rect 30362 921 30542 20454
rect 26498 880 26678 881
rect 30357 743 30363 921
rect 30541 743 30547 921
rect 30362 742 30542 743
<< via3 >>
rect 21588 39454 21652 39518
rect 23244 38460 23308 38524
rect 22140 38038 22204 38102
rect 22692 38092 22756 38156
rect 220 19758 574 20124
rect 3099 17643 3497 18041
rect 26499 881 26677 1059
rect 30363 743 30541 921
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 200 20124 600 44152
rect 200 19758 220 20124
rect 574 19758 600 20124
rect 200 1000 600 19758
rect 800 18042 1200 44152
rect 21590 39519 21650 45152
rect 21587 39518 21653 39519
rect 21587 39454 21588 39518
rect 21652 39454 21653 39518
rect 21587 39453 21653 39454
rect 22142 38103 22202 45152
rect 22694 38157 22754 45152
rect 23246 38525 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 23243 38524 23309 38525
rect 23243 38460 23244 38524
rect 23308 38460 23309 38524
rect 23243 38459 23309 38460
rect 22691 38156 22757 38157
rect 22139 38102 22205 38103
rect 22139 38038 22140 38102
rect 22204 38038 22205 38102
rect 22691 38092 22692 38156
rect 22756 38092 22757 38156
rect 22691 38091 22757 38092
rect 22139 38037 22205 38038
rect 800 18041 3498 18042
rect 800 17643 3099 18041
rect 3497 17643 3498 18041
rect 800 17642 3498 17643
rect 800 1000 1200 17642
rect 26498 1059 26678 1060
rect 26498 881 26499 1059
rect 26677 881 26678 1059
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 881
rect 30362 921 30542 922
rect 30362 743 30363 921
rect 30541 743 30542 921
rect 30362 0 30542 743
use alt  alt_0
timestamp 1762226203
transform 1 0 18204 0 1 19994
box -3708 -3142 4491 1400
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
