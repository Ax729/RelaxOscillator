magic
tech sky130A
magscale 1 2
timestamp 1760057311
<< nwell >>
rect -7886 4218 -7824 4256
rect -7624 4116 -7568 4144
<< pdiff >>
rect -7825 4218 -7824 4256
<< poly >>
rect -7852 4040 -7796 4050
<< locali >>
rect -7624 4116 -7568 4144
rect -7852 4040 -7798 4050
rect -6149 3358 -6085 3364
rect -6149 3262 -6085 3272
<< viali >>
rect -6119 1990 -6055 2054
<< metal1 >>
rect -8992 4828 -4894 4830
rect -8992 4826 -4134 4828
rect -8992 4726 -4070 4826
rect -8992 4596 -8904 4726
rect -4896 4724 -4070 4726
rect -4150 4720 -4070 4724
rect -8992 4490 -8902 4596
rect -8990 4086 -8902 4490
rect -7320 4342 -6764 4390
rect -7870 4116 -7110 4144
rect -9404 4076 -8576 4086
rect -7870 4078 -7836 4116
rect -7160 4078 -7110 4116
rect -9404 4038 -8086 4076
rect -7980 4058 -7110 4078
rect -7980 4038 -7108 4058
rect -8990 3344 -8902 4038
rect -8642 4028 -8086 4038
rect -7172 3652 -7108 4038
rect -6902 3652 -6832 4342
rect -4150 4041 -4074 4720
rect -4150 4040 -4073 4041
rect -4160 3964 -4150 4040
rect -4074 3964 -4064 4040
rect -7324 3598 -6832 3652
rect -7324 3578 -6878 3598
rect -6150 3584 -5700 3630
rect -7172 3346 -7108 3578
rect -4150 3534 -4073 3964
rect -8990 3340 -8572 3344
rect -7178 3340 -7102 3346
rect -8990 3336 -8396 3340
rect -7970 3338 -7172 3340
rect -8346 3336 -7172 3338
rect -8990 3306 -7172 3336
rect -8990 3304 -8902 3306
rect -8796 3302 -7172 3306
rect -8596 3300 -7172 3302
rect -8596 3298 -8196 3300
rect -7288 3060 -7172 3106
rect -8296 2578 -8250 2878
rect -8296 2542 -7922 2578
rect -8848 2038 -8062 2040
rect -9090 1998 -8062 2038
rect -7966 2004 -7930 2542
rect -7328 2304 -7172 2340
rect -7680 2030 -7592 2032
rect -7680 2002 -7172 2030
rect -7600 2000 -7172 2002
rect -7108 3300 -6714 3340
rect -4149 3330 -4073 3534
rect -6092 3308 -5588 3326
rect -6130 3280 -5588 3308
rect -4150 3300 -4072 3330
rect -2534 3302 -2028 3304
rect -4278 3260 -3646 3300
rect -3028 3212 -2028 3302
rect -3028 3210 -2522 3212
rect -7108 3060 -6850 3106
rect -6136 3052 -5698 3096
rect -4294 3020 -3830 3084
rect -6070 2354 -5560 2408
rect -4272 2380 -3768 2426
rect -7108 2304 -6814 2340
rect -2926 2134 -2428 2136
rect -6125 2054 -6049 2066
rect -5882 2054 -4360 2112
rect -4014 2098 -3690 2128
rect -4234 2096 -3690 2098
rect -4234 2066 -3910 2096
rect -2926 2062 -1992 2134
rect -2490 2060 -1992 2062
rect -7038 2030 -6682 2042
rect -7108 2012 -6682 2030
rect -7108 2000 -6898 2012
rect -9090 1996 -8520 1998
rect -9090 1862 -9004 1996
rect -6125 1990 -6119 2054
rect -6055 2048 -4360 2054
rect -6055 1990 -5818 2048
rect -6125 1978 -6049 1990
rect -4248 1862 -3744 1908
rect -9092 1816 -9004 1862
rect -9092 1536 -9006 1816
rect -6086 1804 -5576 1858
rect -7320 1748 -6810 1802
rect -9094 1386 -9006 1536
rect -7338 1486 -6952 1550
rect -9094 1246 -9008 1386
rect -9094 1244 -8042 1246
rect -9248 1202 -8042 1244
rect -7966 1244 -7894 1248
rect -7966 1242 -7858 1244
rect -7774 1242 -7050 1246
rect -9248 1198 -9008 1202
rect -7966 1200 -7050 1242
rect -9094 628 -9008 1198
rect -7898 1196 -7050 1200
rect -7826 1194 -7050 1196
rect -7766 988 -7712 1194
rect -7772 942 -7718 976
rect -7762 906 -7708 942
rect -7762 904 -7194 906
rect -7150 904 -7050 1194
rect -7762 838 -7046 904
rect -7240 836 -7046 838
rect -9094 626 -4916 628
rect -9094 622 -4476 626
rect -9094 536 -3912 622
rect -4936 534 -3912 536
rect -4498 530 -3912 534
<< via1 >>
rect -4150 3964 -4074 4040
rect -7172 2000 -7108 3340
<< metal2 >>
rect -4150 4040 -4074 4050
rect -4150 3954 -4074 3964
rect -7310 3842 -7012 3846
rect -7310 3794 -7004 3842
rect -8628 3340 -8070 3346
rect -8954 3338 -8070 3340
rect -8958 3306 -8070 3338
rect -7172 3340 -7108 3346
rect -8958 3300 -8396 3306
rect -8958 2878 -8880 3300
rect -8958 2842 -8258 2878
rect -7968 2648 -7924 3334
rect -9004 2644 -8724 2646
rect -9004 2642 -8452 2644
rect -8244 2642 -7918 2648
rect -9004 2618 -7918 2642
rect -9002 2614 -8192 2618
rect -7968 2616 -7924 2618
rect -9002 2468 -8914 2614
rect -8472 2612 -8192 2614
rect -9002 2404 -8912 2468
rect -9000 2040 -8912 2404
rect -9000 2036 -8900 2040
rect -9000 2030 -8516 2036
rect -8080 2032 -7478 2036
rect -8314 2030 -7478 2032
rect -9000 2002 -7478 2030
rect -8950 2000 -7478 2002
rect -7054 3092 -7004 3794
rect -4316 3542 -3848 3628
rect -4568 3306 -4088 3308
rect -4952 3270 -4088 3306
rect -4952 3268 -4070 3270
rect -4952 3266 -4408 3268
rect -7054 3046 -6828 3092
rect -4144 2868 -4070 3268
rect -5922 2574 -4966 2580
rect -5922 2536 -4188 2574
rect -8638 1996 -7916 2000
rect -8638 1994 -8240 1996
rect -7172 1196 -7108 2000
rect -7054 2316 -6850 2348
rect -7054 1496 -6966 2316
rect -5920 2112 -5874 2536
rect -5144 2530 -4188 2536
rect -4242 2528 -4194 2530
rect -5920 2110 -5318 2112
rect -5920 2076 -4972 2110
rect -5570 2074 -4972 2076
rect -4260 2098 -4222 2182
rect -4136 2098 -4090 2868
rect -4260 2088 -4090 2098
rect -4260 2066 -4092 2088
rect -4014 1888 -3910 2084
rect -6864 1004 -6792 1820
rect -4016 1712 -3910 1888
rect -4018 1662 -3910 1712
rect -4018 1356 -3912 1662
rect -7328 950 -6792 1004
rect -6864 948 -6792 950
rect -4022 1330 -3912 1356
rect -4022 608 -3916 1330
<< metal3 >>
rect -4242 3300 -4182 3322
rect -4242 3260 -4180 3300
rect -4240 2590 -4180 3260
rect -4240 2528 -4174 2590
use sky130_fd_sc_hd__nand2_8  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -8744 0 1 3824
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x2
timestamp 1704896540
transform 1 0 -8732 0 1 3086
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x3
timestamp 1704896540
transform 1 0 -8732 0 1 1780
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x4
timestamp 1704896540
transform 1 0 -8716 0 1 986
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -6896 0 1 3076
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x6
timestamp 1704896540
transform 1 0 -6866 0 1 1796
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -5710 0 1 3052
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  x8
timestamp 1704896540
transform 1 0 -5668 0 1 1860
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -3888 0 1 3046
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x10
timestamp 1704896540
transform 1 0 -3784 0 1 1882
box -38 -48 1142 592
<< end >>
